toto * tutu;
