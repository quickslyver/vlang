package toto is

 function f(a,b:integer)return integer --test function
 is
   return a+b;
 end function;
end package toto;

